-- PWM_Lkup.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PWM_Lkup is
	port (
		addr       : in  std_logic_vector(8 downto 0)  := (others => '0'); --       addr.addr
		data_valid : out std_logic;                                        -- data_valid.data_valid
		dataout    : out std_logic_vector(15 downto 0);                    --    dataout.dataout
		nbusy      : out std_logic;                                        --      nbusy.nbusy
		nread      : in  std_logic                     := '0'              --      nread.nread
	);
end entity PWM_Lkup;

architecture rtl of PWM_Lkup is
	component PWM_Lkup_ufm_parallel_0 is
		port (
			addr       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- addr
			nread      : in  std_logic                     := 'X';             -- nread
			dataout    : out std_logic_vector(15 downto 0);                    -- dataout
			nbusy      : out std_logic;                                        -- nbusy
			data_valid : out std_logic                                         -- data_valid
		);
	end component PWM_Lkup_ufm_parallel_0;

begin

	ufm_parallel_0 : component PWM_Lkup_ufm_parallel_0
		port map (
			addr       => addr,       --       addr.addr
			nread      => nread,      --      nread.nread
			dataout    => dataout,    --    dataout.dataout
			nbusy      => nbusy,      --      nbusy.nbusy
			data_valid => data_valid  -- data_valid.data_valid
		);

end architecture rtl; -- of PWM_Lkup
